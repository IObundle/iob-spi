`define SPI_ADDR_W 3 // data_width
`define SPI_DATA_W 32 // data_width


// MEMORY MAP
`define SPI_INTRRPT_EN 0
`define SPI_READY 1
`define SPI_TX 2
`define SPI_RX 3
`define DUMMY_REG 7
