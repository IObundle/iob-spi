`define SPI_ADDR_W 2 // data_width
`define SPI_DATA_W 32 // data_width


// MEMORY MAP

`define SPI_START 0
`define SPI_READY 1
`define SPI_TX 2
`define SPI_RX 3
