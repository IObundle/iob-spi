`define	FL_ADDR_W	4	
`define	FL_WDATA_W	32	
`ifndef
	`define	DATA_W	32
`endif
